//Including all the files in the design
//This is the integration file

`include "Shift_Unit.v"  //done
`include "ALU.v"         //done
`include "Misc.v"        //done
`include "Multiplexers.v" //done
`include "Register_Bank.v"  //done
`include "Data_memory.v"   //done
`include "moore_control_unit.v"  //done
`include "IFstage.v"  //done


// Integrating hardware to build Datapath

module processor_datapath(output [3:0] out_15_12,output isZero/*(Zeroflag)*/,
input clk,input IR_write,input PCwritefinal,/*(Final PC Control signal including BE,BNE,Zeroflag)*/input RegDst,input RegWrite,
input MemtoReg,input MDRwrite/*(Control signal enabling write into MDR)*/,input ALUoutwrite/*(Control signal enabling write into ALUOut)*/,
input [1:0] ALUop,input [1:0] ALUSrcA,input [2:0] ALUSrcB,input Shift,input [1:0] PCsrc,
input MemRead,input MemWrite,input reset); //the control signals not specified in comments either have the usual meaning or specified seperately control unit
wire [15:0] PCin;
wire [15:0] Instruction; 
wire [15:0] PCout;
wire [15:0] PCout1; //PC was declared as two units. One used as a data holding unit, the other performing normal function as a PC does.
wire [3:0] out_11_8; //Instruction[11:8]
wire [3:0] out_7_4;  //Instruction[7:4]
wire [3:0] out_3_0;  //Instruction[3:0]
wire [3:0] Write_register; //Destination Register
wire [3:0] Append11_out; 
wire [3:0] Append10_out;
wire [15:0] Write_data;
wire [15:0] A;           // A,B,C,D,E act as intermediate registers between Register Bank and ALU
wire [15:0] B;  
wire [15:0] C;
wire [15:0] D;
wire [15:0] E;
wire [15:0] ALUout;
wire [15:0] mdr_in;
wire [15:0] mdr_out;
wire [15:0] mux_B_2; //inputs of multiplexer feeding to ALUinB
wire [15:0] mux_B_1; //inputs of multiplexer feeding to ALUinB
wire [15:0] mux_B_4; //inputs of multiplexer feeding to ALUinB
wire [15:0] mux_B_3; //inputs of multiplexer feeding to ALUinB
wire [15:0] mux_B_0; //inputs of multiplexer feeding to ALUinB
wire [15:0] ALUinA; //inputs of ALU
wire [15:0] ALUinB; //inputs of ALU
wire [15:0] ALUout1; //output of ALU, input of ALUout
wire [15:0] Shiftout; //Output of Shifting unit created
wire [15:0] result;   //Output of Shift Multiplexer i.e if(Shift instruction)=> result= o/p of Shift Unit; else result=>ALUout


PC_latch IF_latch( PCin,PCwritefinal,reset,PCout1);  //Instantiating all the modules pertinent to the design (names of the modules speak for themselves)
PC_reg IF_reg(clk,PCout1,PCout);
Instruction_memory IM(PCout,Instruction);
IR Instruction_register(Instruction,IR_write,out_15_12,out_11_8,out_7_4,out_3_0);

append_11 append11_mod({out_15_12,out_11_8,out_7_4,out_3_0},Append11_out); //append 10,11 are taken from load/store instructions.
append_10 append10_mod({out_15_12,out_11_8,out_7_4,out_3_0},Append10_out);

Register_Bank Reg_Bank(RegWrite,out_11_8,out_7_4,out_3_0,Append10_out,Append11_out,Write_register,Write_data,clk,A,B,C,D,E);

sign_extend_8bits se_8({out_7_4,out_3_0},mux_B_2);
zeros_extend ze_8({out_7_4,out_3_0},mux_B_1);
left_shift_sign_extend lsse({8'd0,out_7_4,out_3_0},mux_B_4);
pad0_sign_extend pse({8'd0,out_7_4,out_3_0},mux_B_3);
sign_extend_12bits se_12({4'd0,out_11_8,out_7_4,out_3_0},mux_B_0);
mux_reg_dst reg_dst_mux(out_11_8,Append11_out,RegDst,Write_register);

mux_4to1_ALU_in1 ALU_A_mux(E,A,C,PCout,ALUSrcA,ALUinA);
mux_8to1_ALU_in2 ALU_B_mux(mux_B_0,mux_B_1,mux_B_2,mux_B_3,mux_B_4,B,ALUinB,ALUSrcB);
memtoreg_mux mem_to_reg(mdr_out,ALUout,MemtoReg,Write_data);

ALU_16bit ALU(ALUinA,ALUinB,ALUop,ALUout1,isZero);
shift_unit SU(C,out_3_0,out_7_4,Shiftout);
shift_mux selector(ALUout1,Shiftout,Shift,result);
ALU_Out result_reg(ALUout,result,ALUoutwrite);
mux_PC_src Address_mux(ALUout,ALUout1,C,PCsrc,PCin);
Data_memory mem(MemRead,MemWrite,ALUout,D,mdr_in); 
mdr_latch MDR(mdr_in,mdr_out,MDRwrite);
endmodule

module PROCESSOR_RISCY_Mark_V(input clk,input reset); //asynchrounous reset given to the processor as an input
wire PCwritefinal,MemtoReg,IRWrite,MemRead,MemWrite,RegWrite,Shift,RegDst,MDRwrite,ALUoutwrite;
wire [1:0] ALUop;
wire [1:0] ALUSrcA;
wire [1:0] PCsrc;
wire [2:0] ALUSrcB;
wire [3:0] OPCODE;
wire isZero;

processor_datapath RISCY_Mark_V_data(OPCODE,isZero,clk,IRWrite,PCwritefinal,
RegDst,RegWrite,MemtoReg,MDRwrite,ALUoutwrite,ALUop,ALUSrcA,ALUSrcB,Shift,
PCsrc,MemRead,MemWrite,reset);                          //instantiation of datapath of processor

processor_control_unit_moore_fsm RISCY_Mark_V_control(PCwritefinal,ALUop,ALUSrcA,
ALUSrcB,MemtoReg,MDRwrite,ALUoutwrite,IRWrite,MemRead,MemWrite,RegWrite,Shift,PCsrc,
RegDst,OPCODE,clk,isZero);                              //instantion of control unit of processor

always @(reset) begin
    if(reset == 1'b1) begin      // Specifying what reset signal does to the register bank
    RISCY_Mark_V_data.Reg_Bank.R0 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R1 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R2 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R3 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R4 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R5 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R6 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R7 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R8 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R9 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R10 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R11 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R12 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R13 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R14 = 16'd0;
    RISCY_Mark_V_data.Reg_Bank.R15 = 16'd0;
    end
    //else if(reset == 1'b0) PCwrite_reg = PCWrite;
end

endmodule

module testbench_abcd();   //test bench for the processor
reg clk;
reg reset;
PROCESSOR_RISCY_Mark_V uut(clk,reset);
initial begin
        clk = 1'b0;
        forever begin
            #2 clk = ~clk;   //clk cycle of 4sec
        end
end
initial begin
    //$dumpfile("testbench_processor.vcd"); //to be used for iverilog users
    //$dumpvars(0,testbench);
    //#10 $display($time,"IF State = %b, PC = %h, PC+2 = %h, Instruction = %h, PCWrite = %h",uut.RISCY_Mark_V_control.present_state,uut.RISCY_Mark_V_data.Address,uut.RISCY_Mark_V_data.ALUout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal);
    reset = 1'b1; 
    #1 reset = 1'b0;  //reset signal active for 1 sec, for initialization of relevant control signals and registers.
    //$monitor($time," uut.RISCY_Mark_V_data.mem.storage[33] = %h , uut.RISCY_Mark_V_data.mem.storage[34] = %h",uut.RISCY_Mark_V_data.mem.storage[33],uut.RISCY_Mark_V_data.mem.storage[34]);
    #2 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);   
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUsrcA=%h ALUsrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  Mem:Address =%h MDR =%h MemRead =%h MemWrite = %h ",uut.RISCY_Mark_V_data.ALUout , uut.RISCY_Mark_V_data.mdr_in ,  uut.RISCY_Mark_V_data.MemRead , uut.RISCY_Mark_V_data.MemWrite);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  Mem:Address =%h Datain =%h MemRead =%h MemWrite = %h ",uut.RISCY_Mark_V_data.ALUout , uut.RISCY_Mark_V_data.D ,  uut.RISCY_Mark_V_data.MemRead , uut.RISCY_Mark_V_data.MemWrite);    
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);       
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);           
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite,uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);       
    #4 $strobe ("  EX :PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);        
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
    
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);   
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h ",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  Mem:Address =%h MDR =%h MemRead =%h MemWrite = %h ",uut.RISCY_Mark_V_data.ALUout , uut.RISCY_Mark_V_data.mdr_in ,  uut.RISCY_Mark_V_data.MemRead , uut.RISCY_Mark_V_data.MemWrite);
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);
    #4 $strobe ("  Mem:Address =%h Datain =%h MemRead =%h MemWrite = %h ",uut.RISCY_Mark_V_data.ALUout , uut.RISCY_Mark_V_data.D ,  uut.RISCY_Mark_V_data.MemRead , uut.RISCY_Mark_V_data.MemWrite);    
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite); 
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);   
    #4 $strobe ("  WB :R0 =%h R1 = %h R2 =%h R3 = %h R4 =%h R5 = %h R6 =%h R7 = %h R8 =%h R9 = %h R10 =%h R11 = %h R12 =%h R13 = %h R14 =%h R15 = %h MemtoReg=%h RegDst=%h RegWrite =%h", uut.RISCY_Mark_V_data.Reg_Bank.R0,uut.RISCY_Mark_V_data.Reg_Bank.R1 ,uut.RISCY_Mark_V_data.Reg_Bank.R2 ,uut.RISCY_Mark_V_data.Reg_Bank.R3 , uut.RISCY_Mark_V_data.Reg_Bank.R4,uut.RISCY_Mark_V_data.Reg_Bank.R5,uut.RISCY_Mark_V_data.Reg_Bank.R6,uut.RISCY_Mark_V_data.Reg_Bank.R7,uut.RISCY_Mark_V_data.Reg_Bank.R8,uut.RISCY_Mark_V_data.Reg_Bank.R9,uut.RISCY_Mark_V_data.Reg_Bank.R10,uut.RISCY_Mark_V_data.Reg_Bank.R11,uut.RISCY_Mark_V_data.Reg_Bank.R12,uut.RISCY_Mark_V_data.Reg_Bank.R13,uut.RISCY_Mark_V_data.Reg_Bank.R14,uut.RISCY_Mark_V_data.Reg_Bank.R15,uut.RISCY_Mark_V_data.MemtoReg,uut.RISCY_Mark_V_data.RegDst,uut.RISCY_Mark_V_data.RegWrite);   
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);       
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);           
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h ALUout=%h ALUinA =%h ALUinB =%h ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite,uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop);       
    #4 $strobe ("  EX :PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);        
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
    #4 $strobe ("  IF: PC=%h Updated PC=%h Instruction=%h PCwritefinal =%h IRwrite =%h ",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.PCout1,uut.RISCY_Mark_V_data.Instruction,uut.RISCY_Mark_V_data.PCwritefinal,uut.RISCY_Mark_V_data.IR_write);
    #4 $strobe ("  ID :PC=%h A=%h B=%h C=%h D=%h E=%h Regwrite=%h",uut.RISCY_Mark_V_data.PCout,uut.RISCY_Mark_V_data.A,uut.RISCY_Mark_V_data.B,uut.RISCY_Mark_V_data.C,uut.RISCY_Mark_V_data.D,uut.RISCY_Mark_V_data.E,uut.RISCY_Mark_V_data.RegWrite);       
    #4 $strobe ("  EX :ALUout=%h ALUinA =%h ALUinB =%H ALUSrcA=%h ALUSrcB=%h  Shift=%h  ALUoutWrite =%h ALUop =%h PCSrc= %h PC=%h",uut.RISCY_Mark_V_data.ALUout,uut.RISCY_Mark_V_data.ALUinA,uut.RISCY_Mark_V_data.ALUinB,uut.RISCY_Mark_V_data.ALUSrcA,uut.RISCY_Mark_V_data.ALUSrcB,uut.RISCY_Mark_V_data.Shift,uut.RISCY_Mark_V_data.ALUoutwrite,uut.RISCY_Mark_V_data.ALUop,uut.RISCY_Mark_V_data.PCsrc,uut.RISCY_Mark_V_data.PCout1);          
      
        //#1000 $finish;
end

endmodule


